-- ----------------------------------------------------------------------------
-- Module:          uzed_top.vhd
-- Description:     Top level module of 6502 based single board computer for
--                  Avnet Microzed 7010 or 7020
-- Author:          George Castillo
-- Date:            20 November 2023
--
-- TODO Supports:
--   - Directive selecting whether to target a Microzed 7010 or 7020 as well
--     as the carrier board to use (if any).
--   - Alternate clock sources to specify
--
-- ----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity uzed_top is
    port (
        DDR_addr            : inout std_logic_vector (14 downto 0);
        DDR_ba              : inout std_logic_vector (2 downto 0);
        DDR_cas_n           : inout std_logic;
        DDR_ck_n            : inout std_logic;
        DDR_ck_p            : inout std_logic;
        DDR_cke             : inout std_logic;
        DDR_cs_n            : inout std_logic;
        DDR_dm              : inout std_logic_vector (3 downto 0);
        DDR_dq              : inout std_logic_vector (31 downto 0);
        DDR_dqs_n           : inout std_logic_vector (3 downto 0);
        DDR_dqs_p           : inout std_logic_vector (3 downto 0);
        DDR_odt             : inout std_logic;
        DDR_ras_n           : inout std_logic;
        DDR_reset_n         : inout std_logic;
        DDR_we_n            : inout std_logic;

        FIXED_IO_ddr_vrn    : inout std_logic;
        FIXED_IO_ddr_vrp    : inout std_logic;
        FIXED_IO_mio        : inout std_logic_vector (53 downto 0);
        FIXED_IO_ps_clk     : inout std_logic;
        FIXED_IO_ps_porb    : inout std_logic;
        FIXED_IO_ps_srstb   : inout std_logic
      );

end entity uzed_top;

architecture structural of uzed_top is

    -- PS7 block design signals. These should be pulled directly from the VHDL wrapper that was
    -- generated by Vivado. Some rearrangement is allowed to logically group related signals but
    -- port widths and names should be untouched.

    -- SBC clock and reset. Much of the SBC logic needs to be run from a 100MHz clock, particularly
    -- the clock and reset generator.
    signal SBC_CLK              : std_logic;
    signal SBC_RSTN             : std_logic;

    -- AXI interface to SBC control and registers
    signal SBC_CTRL_araddr      : std_logic_vector(31 downto 0);
    signal SBC_CTRL_arburst     : std_logic_vector(1 downto 0);
    signal SBC_CTRL_arcache     : std_logic_vector(3 downto 0);
    signal SBC_CTRL_arid        : std_logic_vector(11 downto 0);
    signal SBC_CTRL_arlen       : std_logic_vector(7 downto 0);
    signal SBC_CTRL_arlock      : std_logic_vector(0 to 0);
    signal SBC_CTRL_arprot      : std_logic_vector(2 downto 0);
    signal SBC_CTRL_arqos       : std_logic_vector(3 downto 0);
    signal SBC_CTRL_arready     : std_logic_vector(0 to 0);
    signal SBC_CTRL_arregion    : std_logic_vector(3 downto 0);
    signal SBC_CTRL_arsize      : std_logic_vector(2 downto 0);
    signal SBC_CTRL_arvalid     : std_logic_vector(0 to 0);
    signal SBC_CTRL_awaddr      : std_logic_vector(31 downto 0);
    signal SBC_CTRL_awburst     : std_logic_vector(1 downto 0);
    signal SBC_CTRL_awcache     : std_logic_vector(3 downto 0);
    signal SBC_CTRL_awid        : std_logic_vector(11 downto 0);
    signal SBC_CTRL_awlen       : std_logic_vector(7 downto 0);
    signal SBC_CTRL_awlock      : std_logic_vector(0 to 0);
    signal SBC_CTRL_awprot      : std_logic_vector(2 downto 0);
    signal SBC_CTRL_awqos       : std_logic_vector(3 downto 0);
    signal SBC_CTRL_awready     : std_logic_vector(0 to 0);
    signal SBC_CTRL_awregion    : std_logic_vector(3 downto 0);
    signal SBC_CTRL_awsize      : std_logic_vector(2 downto 0);
    signal SBC_CTRL_awvalid     : std_logic_vector(0 to 0);
    signal SBC_CTRL_bid         : std_logic_vector(11 downto 0);
    signal SBC_CTRL_bready      : std_logic_vector(0 to 0);
    signal SBC_CTRL_bresp       : std_logic_vector(1 downto 0);
    signal SBC_CTRL_bvalid      : std_logic_vector(0 to 0);
    signal SBC_CTRL_rdata       : std_logic_vector(31 downto 0);
    signal SBC_CTRL_rid         : std_logic_vector(11 downto 0);
    signal SBC_CTRL_rlast       : std_logic_vector(0 to 0);
    signal SBC_CTRL_rready      : std_logic_vector(0 to 0);
    signal SBC_CTRL_rresp       : std_logic_vector(1 downto 0);
    signal SBC_CTRL_rvalid      : std_logic_vector(0 to 0);
    signal SBC_CTRL_wdata       : std_logic_vector(31 downto 0);
    signal SBC_CTRL_wlast       : std_logic_vector(0 to 0);
    signal SBC_CTRL_wready      : std_logic_vector(0 to 0);
    signal SBC_CTRL_wstrb       : std_logic_vector(3 downto 0);
    signal SBC_CTRL_wvalid      : std_logic_vector(0 to 0);

    -- AXI to block RAM interface for EEPROM emulator
    signal SBC_EEPROM_addr      : std_logic_vector(12 downto 0);
    signal SBC_EEPROM_clk       : std_logic;
    signal SBC_EEPROM_din       : std_logic_vector(31 downto 0);
    signal SBC_EEPROM_dout      : std_logic_vector(31 downto 0);
    signal SBC_EEPROM_en        : std_logic;
    signal SBC_EEPROM_rst       : std_logic;
    signal SBC_EEPROM_we        : std_logic_vector(3 downto 0);

    -- AXI to block RAM interface for SRAM emulator
    signal SBC_SRAM_addr        : std_logic_vector(12 downto 0);
    signal SBC_SRAM_clk         : std_logic;
    signal SBC_SRAM_din         : std_logic_vector(31 downto 0);
    signal SBC_SRAM_dout        : std_logic_vector(31 downto 0);
    signal SBC_SRAM_en          : std_logic;
    signal SBC_SRAM_rst         : std_logic;
    signal SBC_SRAM_we          : std_logic_vector(3 downto 0);

    -- Hardware timers (TTC0)
    signal TTC0_WAVE0           : std_logic;
    signal TTC0_WAVE1           : std_logic;
    signal TTC0_WAVE2           : std_logic;

begin

    -- Instantiates the Zynq PS block design with exported AXI interfaces, clocks, resets, block RAM
    -- interfaces, and all other supporting signals. In general, this should be wired up as is with
    -- port names as signals (so that macros can easily process it if changes are necessary) and
    -- then signals routed to the appropriate locations, or as top level port names (e.g., DDR and
    -- FIXED_IO signals).
    ps7_bd: entity work.ps7_wrapper
    port map (
        DDR_addr            => DDR_addr,            -- STD_LOGIC_VECTOR ( 14 downto 0 )
        DDR_ba              => DDR_ba,              -- STD_LOGIC_VECTOR ( 2 downto 0 )
        DDR_cas_n           => DDR_cas_n,           -- STD_LOGIC
        DDR_ck_n            => DDR_ck_n,            -- STD_LOGIC
        DDR_ck_p            => DDR_ck_p,            -- STD_LOGIC
        DDR_cke             => DDR_cke,             -- STD_LOGIC
        DDR_cs_n            => DDR_cs_n,            -- STD_LOGIC
        DDR_dm              => DDR_dm,              -- STD_LOGIC_VECTOR ( 3 downto 0 )
        DDR_dq              => DDR_dq,              -- STD_LOGIC_VECTOR ( 31 downto 0 )
        DDR_dqs_n           => DDR_dqs_n,           -- STD_LOGIC_VECTOR ( 3 downto 0 )
        DDR_dqs_p           => DDR_dqs_p,           -- STD_LOGIC_VECTOR ( 3 downto 0 )
        DDR_odt             => DDR_odt,             -- STD_LOGIC
        DDR_ras_n           => DDR_ras_n,           -- STD_LOGIC
        DDR_reset_n         => DDR_reset_n,         -- STD_LOGIC
        DDR_we_n            => DDR_we_n,            -- STD_LOGIC
        FIXED_IO_ddr_vrn    => FIXED_IO_ddr_vrn,    -- STD_LOGIC
        FIXED_IO_ddr_vrp    => FIXED_IO_ddr_vrp,    -- STD_LOGIC
        FIXED_IO_mio        => FIXED_IO_mio,        -- STD_LOGIC_VECTOR ( 53 downto 0 )
        FIXED_IO_ps_clk     => FIXED_IO_ps_clk,     -- STD_LOGIC
        FIXED_IO_ps_porb    => FIXED_IO_ps_porb,    -- STD_LOGIC
        FIXED_IO_ps_srstb   => FIXED_IO_ps_srstb,   -- STD_LOGIC
        SBC_CLK             => SBC_CLK,             -- STD_LOGIC
        SBC_CTRL_araddr     => SBC_CTRL_araddr,     -- STD_LOGIC_VECTOR ( 31 downto 0 )
        SBC_CTRL_arburst    => SBC_CTRL_arburst,    -- STD_LOGIC_VECTOR ( 1 downto 0 )
        SBC_CTRL_arcache    => SBC_CTRL_arcache,    -- STD_LOGIC_VECTOR ( 3 downto 0 )
        SBC_CTRL_arid       => SBC_CTRL_arid,       -- STD_LOGIC_VECTOR ( 11 downto 0 )
        SBC_CTRL_arlen      => SBC_CTRL_arlen,      -- STD_LOGIC_VECTOR ( 7 downto 0 )
        SBC_CTRL_arlock     => SBC_CTRL_arlock,     -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_arprot     => SBC_CTRL_arprot,     -- STD_LOGIC_VECTOR ( 2 downto 0 )
        SBC_CTRL_arqos      => SBC_CTRL_arqos,      -- STD_LOGIC_VECTOR ( 3 downto 0 )
        SBC_CTRL_arready    => SBC_CTRL_arready,    -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_arregion   => SBC_CTRL_arregion,   -- STD_LOGIC_VECTOR ( 3 downto 0 )
        SBC_CTRL_arsize     => SBC_CTRL_arsize,     -- STD_LOGIC_VECTOR ( 2 downto 0 )
        SBC_CTRL_arvalid    => SBC_CTRL_arvalid,    -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_awaddr     => SBC_CTRL_awaddr,     -- STD_LOGIC_VECTOR ( 31 downto 0 )
        SBC_CTRL_awburst    => SBC_CTRL_awburst,    -- STD_LOGIC_VECTOR ( 1 downto 0 )
        SBC_CTRL_awcache    => SBC_CTRL_awcache,    -- STD_LOGIC_VECTOR ( 3 downto 0 )
        SBC_CTRL_awid       => SBC_CTRL_awid,       -- STD_LOGIC_VECTOR ( 11 downto 0 )
        SBC_CTRL_awlen      => SBC_CTRL_awlen,      -- STD_LOGIC_VECTOR ( 7 downto 0 )
        SBC_CTRL_awlock     => SBC_CTRL_awlock,     -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_awprot     => SBC_CTRL_awprot,     -- STD_LOGIC_VECTOR ( 2 downto 0 )
        SBC_CTRL_awqos      => SBC_CTRL_awqos,      -- STD_LOGIC_VECTOR ( 3 downto 0 )
        SBC_CTRL_awready    => SBC_CTRL_awready,    -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_awregion   => SBC_CTRL_awregion,   -- STD_LOGIC_VECTOR ( 3 downto 0 )
        SBC_CTRL_awsize     => SBC_CTRL_awsize,     -- STD_LOGIC_VECTOR ( 2 downto 0 )
        SBC_CTRL_awvalid    => SBC_CTRL_awvalid,    -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_bid        => SBC_CTRL_bid,        -- STD_LOGIC_VECTOR ( 11 downto 0 )
        SBC_CTRL_bready     => SBC_CTRL_bready,     -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_bresp      => SBC_CTRL_bresp,      -- STD_LOGIC_VECTOR ( 1 downto 0 )
        SBC_CTRL_bvalid     => SBC_CTRL_bvalid,     -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_rdata      => SBC_CTRL_rdata,      -- STD_LOGIC_VECTOR ( 31 downto 0 )
        SBC_CTRL_rid        => SBC_CTRL_rid,        -- STD_LOGIC_VECTOR ( 11 downto 0 )
        SBC_CTRL_rlast      => SBC_CTRL_rlast,      -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_rready     => SBC_CTRL_rready,     -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_rresp      => SBC_CTRL_rresp,      -- STD_LOGIC_VECTOR ( 1 downto 0 )
        SBC_CTRL_rvalid     => SBC_CTRL_rvalid,     -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_wdata      => SBC_CTRL_wdata,      -- STD_LOGIC_VECTOR ( 31 downto 0 )
        SBC_CTRL_wlast      => SBC_CTRL_wlast,      -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_wready     => SBC_CTRL_wready,     -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_CTRL_wstrb      => SBC_CTRL_wstrb,      -- STD_LOGIC_VECTOR ( 3 downto 0 )
        SBC_CTRL_wvalid     => SBC_CTRL_wvalid,     -- STD_LOGIC_VECTOR ( 0 to 0 )
        SBC_EEPROM_addr     => SBC_EEPROM_addr,     -- STD_LOGIC_VECTOR ( 12 downto 0 )
        SBC_EEPROM_clk      => SBC_EEPROM_clk,      -- STD_LOGIC
        SBC_EEPROM_din      => SBC_EEPROM_din,      -- STD_LOGIC_VECTOR ( 31 downto 0 )
        SBC_EEPROM_dout     => SBC_EEPROM_dout,     -- STD_LOGIC_VECTOR ( 31 downto 0 )
        SBC_EEPROM_en       => SBC_EEPROM_en,       -- STD_LOGIC
        SBC_EEPROM_rst      => SBC_EEPROM_rst,      -- STD_LOGIC
        SBC_EEPROM_we       => SBC_EEPROM_we,       -- STD_LOGIC_VECTOR ( 3 downto 0 )
        SBC_RSTN            => SBC_RSTN,            -- STD_LOGIC
        SBC_SRAM_addr       => SBC_SRAM_addr,       -- STD_LOGIC_VECTOR ( 12 downto 0 )
        SBC_SRAM_clk        => SBC_SRAM_clk,        -- STD_LOGIC
        SBC_SRAM_din        => SBC_SRAM_din,        -- STD_LOGIC_VECTOR ( 31 downto 0 )
        SBC_SRAM_dout       => SBC_SRAM_dout,       -- STD_LOGIC_VECTOR ( 31 downto 0 )
        SBC_SRAM_en         => SBC_SRAM_en,         -- STD_LOGIC
        SBC_SRAM_rst        => SBC_SRAM_rst,        -- STD_LOGIC
        SBC_SRAM_we         => SBC_SRAM_we,         -- STD_LOGIC_VECTOR ( 3 downto 0 )
        TTC0_WAVE0          => TTC0_WAVE0,          -- STD_LOGIC
        TTC0_WAVE1          => TTC0_WAVE1,          -- STD_LOGIC
        TTC0_WAVE2          => TTC0_WAVE2           -- STD_LOGIC
    );

    sbc_core_i0: entity work.sbc_core
    generic map (
        VENDOR                  => "XILINX",
        TARGET                  => "7SERIES",
        ADD_CLK_IBUF            => false,
        ADD_RST_IBUF            => false,
        REF_RST_LENGTH          => 8,
        MST_RST_LENGTH          => 8,
        PPU_EN_RST_LENGTH       => 4,
        CPU_EN_RST_LENGTH       => 4
    )
    port map (
        clk_ext                 => SBC_CLK,             -- in    std_logic;
        rst_ext                 => not SBC_RSTN,        -- in    std_logic;
        ext_rom_clk             => SBC_EEPROM_clk,      -- in    std_logic;
        ext_rom_rst             => SBC_EEPROM_rst,      -- in    std_logic;
        ext_rom_en              => SBC_EEPROM_en,       -- in    std_logic;
        ext_rom_we              => SBC_EEPROM_we,       -- in    std_logic_vector(3 downto 0);
        ext_rom_addr            => SBC_EEPROM_addr,     -- in    std_logic_vector(12 downto 0);
        ext_rom_wr_data         => SBC_EEPROM_din,      -- in    std_logic_vector(31 downto 0);
        ext_rom_rd_data         => SBC_EEPROM_dout,     -- out   std_logic_vector(31 downto 0);
        ext_sram_clk            => SBC_SRAM_clk,        -- in    std_logic;
        ext_sram_rst            => SBC_SRAM_rst,        -- in    std_logic;
        ext_sram_en             => SBC_SRAM_en,         -- in    std_logic;
        ext_sram_we             => SBC_SRAM_we,         -- in    std_logic_vector(3 downto 0);
        ext_sram_addr           => SBC_SRAM_addr,       -- in    std_logic_vector(12 downto 0);
        ext_sram_wr_data        => SBC_SRAM_din,        -- in    std_logic_vector(31 downto 0);
        ext_sram_rd_data        => SBC_SRAM_dout        -- out   std_logic_vector(31 downto 0)
    );

end architecture structural;

