-- Clock and reset generation and distribution
--
-- This module receives all four fabric clocks 
-- 
entity clk_rst
    port (
        
